library ieee;
use ieee.std_logic_1164.all;

package constants is
	-- Configuration
	constant WORD_SIZE : natural := 32;

end package constants;

package body constants is
end package body constants;
